`default_nettype none

module dependency_detecter
  (

   input wire clk,
   input wire rstn
  );
endmodule
`default_nettype wire
